* D:\Designs\Pspice\RF_Detector.sch

* Schematics Version 9.2
* Sun Jun 07 21:29:03 2009


.PARAM         in=10m 

** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "RF_Detector.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
