* D:\Designs\Pspice\diodo.sch

* Schematics Version 9.2
* Sun Jun 07 19:28:43 2009


.PARAM         in=0 

** Analysis setup **
.DC LIN PARAM in 0V .7V 10uV 
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "diodo.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
