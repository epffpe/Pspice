* D:\Designs\Pspice\ModuladorAM.sch

* Schematics Version 9.2
* Tue Dec 16 01:39:06 2008



** Analysis setup **
.tran 0ns 50us 1u 1n
.OP 


* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "ModuladorAM.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
