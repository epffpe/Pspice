* D:\Designs\Pspice\DemFMCuadratura.sch

* Schematics Version 9.2
* Wed Jan 07 04:34:41 2009



** Analysis setup **
.tran 0ns 2ms 0.2m 1000n
.OP 


* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "DemFMCuadratura.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
