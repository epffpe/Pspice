* D:\Designs\Pspice\salidaGilbert.sch

* Schematics Version 9.2
* Sun Dec 14 14:17:52 2008



** Analysis setup **
.tran 0ns 20us 0 1n
.OP 


* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "salidaGilbert.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
