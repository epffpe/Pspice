* D:\Designs\Pspice\ClaseC_5V.sch

* Schematics Version 9.2
* Thu Nov 27 23:53:14 2008



** Analysis setup **
.ac LIN 1001 1meg 100meg
.OP 


* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "ClaseC_5V.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
