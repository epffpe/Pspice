* D:\Designs\Pspice\switch.sch

* Schematics Version 9.2
* Sun Dec 14 22:23:23 2008



** Analysis setup **
.tran 0ns 2ms 0 20n
.OP 


* From [PSPICE NETLIST] section of D:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "switch.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
